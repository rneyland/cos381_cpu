library ieee;
use ieee.std_logic_1164.all;

entity Shift32_tb is
end Shift32_tb;

architecture Test of Shift32_tb is
    signal Input, Amount, Output:		std_logic_vector(31 downto 0);
    signal Right, Negative, CarryOut:	std_logic;
begin
    Shift32: entity work.Shift32(rtl) port map (Input, Amount, Right, Output, Negative, CarryOut);
	process
        type PatternType is record
            Input, Amount:		std_logic_vector(31 downto 0);
            Right:				std_logic;
            Output: 			std_logic_vector(31 downto 0);
			Negative, CarryOut:	std_logic;
        end record;
        type PatternArray is array (natural range <>) of PatternType;
        constant Patterns: PatternArray := 
			 -- left shift tests
            (("00000000000000000000000000000001", "00000000000000000000000000000000", '0', "00000000000000000000000000000001", '0', '0'),
			 ("11111111111111111111111111111111", "00000000000000000000000000000000", '0', "11111111111111111111111111111111", '1', '0'),					
			 ("00000000000000000000000000000001", "00000000000000000000000000000001", '0', "00000000000000000000000000000010", '0', '0'),
             ("00000000000000000000000000000001", "00000000000000000000000000000010", '0', "00000000000000000000000000000100", '0', '0'),
             ("00000000000000000000000000000001", "00000000000000000000000000000100", '0', "00000000000000000000000000010000", '0', '0'),
             ("00000000000000000000000000000001", "00000000000000000000000000001000", '0', "00000000000000000000000100000000", '0', '0'),
             ("00000000000000000000000000000001", "00000000000000000000000000010000", '0', "00000000000000010000000000000000", '0', '0'),
             ("00000000000000000000000000000001", "00000000000000000000000000011111", '0', "10000000000000000000000000000000", '1', '0'),
			 ("10000000000000000000000000000000", "00000000000000000000000000000001", '0', "00000000000000000000000000000000", '0', '1'),	
			 ("00100000000000000000000000000000", "00000000000000000000000000000011", '0', "00000000000000000000000000000000", '0', '1'),
			 ("00000000000000000000000000000010", "00000000000000000000000000011111", '0', "00000000000000000000000000000000", '0', '1'),
			 -- right shift tests
			 ("10000000000000000000000000000000", "00000000000000000000000000000000", '1', "10000000000000000000000000000000", '1', '0'),
			 ("11111111111111111111111111111111", "00000000000000000000000000000000", '1', "11111111111111111111111111111111", '1', '0'),	
			 ("10000000000000000000000000000000", "00000000000000000000000000000001", '1', "01000000000000000000000000000000", '0', '0'),
			 ("10000000000000000000000000000000", "00000000000000000000000000000010", '1', "00100000000000000000000000000000", '0', '0'),
			 ("10000000000000000000000000000000", "00000000000000000000000000000100", '1', "00001000000000000000000000000000", '0', '0'),
             ("10000000000000000000000000000000", "00000000000000000000000000001000", '1', "00000000100000000000000000000000", '0', '0'),
             ("10000000000000000000000000000000", "00000000000000000000000000010000", '1', "00000000000000001000000000000000", '0', '0'),
			 ("10000000000000000000000000000000", "00000000000000000000000000011111", '1', "00000000000000000000000000000001", '0', '0'),
			 ("00000000000000000000000000000001", "00000000000000000000000000000001", '1', "00000000000000000000000000000000", '0', '1'),
			 ("00000000000000000000000000000100", "00000000000000000000000000000011", '1', "00000000000000000000000000000000", '0', '1'),
			 ("01000000000000000000000000000000", "00000000000000000000000000011111", '1', "00000000000000000000000000000000", '0', '1'));
	begin
        for i in Patterns'range loop
            Input   <= Patterns(i).Input;
            Amount	<= Patterns(i).Amount;
            Right   <= Patterns(i).Right;
            wait for 1 ns;
            assert Output = Patterns(i).Output
                report "bad Output bits" severity error;
			assert CarryOut = Patterns(i).CarryOut
				report "bad CarryOut bit" severity error;
            assert Negative = Patterns(i).Negative
                report "bad Negative bit" severity error;
        end loop;
        assert false report "end of test" severity note;
        wait;
    end process;
end Test;
